module InstMem(
    input [31:0] address,
    output reg [31:0] inst
);
    
    always @(*)
        case (address[10:2])  // ���512��ָ��
//            9'd0: inst <= 32'h2009000c;
//            9'd1: inst <= 32'h200a0014;
//            9'd2: inst <= 32'h012a4020;
//            9'd3: inst <= 32'h01495822;
//            9'd4: inst <= 32'h200d0010;
//            9'd5: inst <= 32'hac0b0000;
//            9'd6: inst <= 32'h8c0c0000;
//            9'd7: inst <= 32'had8d0000;
//            9'd8: inst <= 32'h200e0014;
//            9'd9: inst <= 32'h114e0000;
//            9'd10: inst <= 32'h000e7080;
//            9'd11: inst <= 32'h0810000a;
9'd0: inst <= 32'h00004020;
9'd1: inst <= 32'h2009003F;
9'd2: inst <= 32'hAD090000;
9'd3: inst <= 32'h21080004;
9'd4: inst <= 32'h20090006;
9'd5: inst <= 32'hAD090000;
9'd6: inst <= 32'h21080004;
9'd7: inst <= 32'h2009005B;
9'd8: inst <= 32'hAD090000;
9'd9: inst <= 32'h21080004;
9'd10: inst <= 32'h2009004F;
9'd11: inst <= 32'hAD090000;
9'd12: inst <= 32'h21080004;
9'd13: inst <= 32'h20090066;
9'd14: inst <= 32'hAD090000;
9'd15: inst <= 32'h21080004;
9'd16: inst <= 32'h2009006D;
9'd17: inst <= 32'hAD090000;
9'd18: inst <= 32'h21080004;
9'd19: inst <= 32'h2009007D;
9'd20: inst <= 32'hAD090000;
9'd21: inst <= 32'h21080004;
9'd22: inst <= 32'h20090007;
9'd23: inst <= 32'hAD090000;
9'd24: inst <= 32'h21080004;
9'd25: inst <= 32'h2009007F;
9'd26: inst <= 32'hAD090000;
9'd27: inst <= 32'h21080004;
9'd28: inst <= 32'h2009006F;
9'd29: inst <= 32'hAD090000;
9'd30: inst <= 32'h21080004;
9'd31: inst <= 32'h200900F7;
9'd32: inst <= 32'hAD090000;
9'd33: inst <= 32'h21080004;
9'd34: inst <= 32'h200900FF;
9'd35: inst <= 32'hAD090000;
9'd36: inst <= 32'h21080004;
9'd37: inst <= 32'h200900B9;
9'd38: inst <= 32'hAD090000;
9'd39: inst <= 32'h21080004;
9'd40: inst <= 32'h200900BF;
9'd41: inst <= 32'hAD090000;
9'd42: inst <= 32'h21080004;
9'd43: inst <= 32'h200900F9;
9'd44: inst <= 32'hAD090000;
9'd45: inst <= 32'h21080004;
9'd46: inst <= 32'h200900F1;
9'd47: inst <= 32'hAD090000;
9'd48: inst <= 32'h21080004;
9'd49: inst <= 32'h0000B820;
9'd50: inst <= 32'h8D110000;
9'd51: inst <= 32'h21050004;
9'd52: inst <= 32'h0C100037;
9'd53: inst <= 32'hAD170000;
9'd54: inst <= 32'h08100059;
9'd55: inst <= 32'h20190001;
9'd56: inst <= 32'h20AB0004;
9'd57: inst <= 32'h02397822;
9'd58: inst <= 32'h19E0001D;
9'd59: inst <= 32'h2338FFFF;
9'd60: inst <= 32'h8D690000;
9'd61: inst <= 32'h216CFFFC;
9'd62: inst <= 32'h07000007;
9'd63: inst <= 32'h22F70001;
9'd64: inst <= 32'h8D8A0000;
9'd65: inst <= 32'h01497822;
9'd66: inst <= 32'h19E00003;
9'd67: inst <= 32'h2318FFFF;
9'd68: inst <= 32'h218CFFFC;
9'd69: inst <= 32'h0810003E;
9'd70: inst <= 32'h230D0001;
9'd71: inst <= 32'h218E0004;
9'd72: inst <= 32'h2338FFFF;
9'd73: inst <= 32'h8D690000;
9'd74: inst <= 32'h216CFFFC;
9'd75: inst <= 32'h030D7822;
9'd76: inst <= 32'h05E00005;
9'd77: inst <= 32'h8D8A0000;
9'd78: inst <= 32'hAD8A0004;
9'd79: inst <= 32'h2318FFFF;
9'd80: inst <= 32'h218CFFFC;
9'd81: inst <= 32'h0810004B;
9'd82: inst <= 32'hADC90000;
9'd83: inst <= 32'h23390001;
9'd84: inst <= 32'h216B0004;
9'd85: inst <= 32'h03317822;
9'd86: inst <= 32'h05E0FFE2;
9'd87: inst <= 32'h08100058;
9'd88: inst <= 32'h03E00008;
9'd89: inst <= 32'h22300001;
9'd90: inst <= 32'h3C014000;
9'd91: inst <= 32'h34210010;
9'd92: inst <= 32'h00018820;
9'd93: inst <= 32'h2009003C;
9'd94: inst <= 32'h12000028;
9'd95: inst <= 32'h21290004;
9'd96: inst <= 32'h8D2A0000;
9'd97: inst <= 32'h2018007D;
9'd98: inst <= 32'h000A5F00;
9'd99: inst <= 32'h000B5F02;
9'd100: inst <= 32'h000B5880;
9'd101: inst <= 32'h8D6F0000;
9'd102: inst <= 32'h21EF0100;
9'd103: inst <= 32'hAE2F0000;
9'd104: inst <= 32'h0C100081;
9'd105: inst <= 32'h000A6600;
9'd106: inst <= 32'h000C6702;
9'd107: inst <= 32'h000C6080;
9'd108: inst <= 32'h8D8F0000;
9'd109: inst <= 32'h21EF0200;
9'd110: inst <= 32'hAE2F0000;
9'd111: inst <= 32'h0C100081;
9'd112: inst <= 32'h000A6D00;
9'd113: inst <= 32'h000D6F02;
9'd114: inst <= 32'h000D6880;
9'd115: inst <= 32'h8DAF0000;
9'd116: inst <= 32'h21EF0400;
9'd117: inst <= 32'hAE2F0000;
9'd118: inst <= 32'h0C100081;
9'd119: inst <= 32'h000A7302;
9'd120: inst <= 32'h000E7080;
9'd121: inst <= 32'h8DCF0000;
9'd122: inst <= 32'h21EF0800;
9'd123: inst <= 32'hAE2F0000;
9'd124: inst <= 32'h0C100081;
9'd125: inst <= 32'h2318FFFF;
9'd126: inst <= 32'h1F00FFE3;
9'd127: inst <= 32'h2210FFFF;
9'd128: inst <= 32'h0810005E;
9'd129: inst <= 32'h3C010000;
9'd130: inst <= 32'h3421C350;
9'd131: inst <= 32'h00014020;
9'd132: inst <= 32'h2108FFFF;
9'd133: inst <= 32'h1D00FFFE;
9'd134: inst <= 32'h03E00008;
9'd135: inst <= 32'hAE200000;
9'd136: inst <= 32'h08100087;




            default: inst <= 32'h0000_0000;
        endcase


endmodule